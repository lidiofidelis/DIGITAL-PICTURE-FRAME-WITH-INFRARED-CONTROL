module ir_encoder(
	input [7:0]data,
	input data_ready,
	input clk,
	output [3:0]controle
);

reg [3:0]temp;

endmodule 